module register(q, d, wrenable, clk);
input d;
input wrenable;
input clk;
output reg q;
always @(posedge clk) begin
	if(wrenable) begin
	q = d;
	end
end
endmodule

module register32(q, d, wrenable, clk);
input[31:0] d;
input wrenable;
input clk;
output reg[31:0] q;

always @(posedge clk) begin
	if(wrenable) begin
	q = d;
	end
end
endmodule

module register32zero(q, d, wrenable, clk);
input[31:0] d;
input wrenable;
input clk;
output reg[31:0] q;
wire zeroenable;

and and1(zeroenable, wrenable, 0);

always @(posedge clk) begin
	if(wrenable) begin
	q = d;
	end
end
endmodule

module mux32to1by1(out, address, inputs);
input[31:0] inputs;
input[4:0] address;
output out;
assign out = inputs[address];
endmodule

module mux32to1by32(out, address, inputs);
//module mux32to1by32(out, address, input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15, input16, input17, input18, input19, input20, input21, input22, input23, input24, input25, input26, input27, input28, input29, input30, input31);
//input[31:0] input0, input1, input2, input3, input4, input5, input6, input7, input8, input9, input10, input11, input12, input13, input14, input15, input16, input17, input18, input19, input20, input21, input22, input23, input24, input25, input26, input27, input28, input29, input30, input31;
input[31:0] inputs[31:0]
input[4:0] address;
output[31:0] out;
wire[31:0] mux[31:0]; // Creates a 2d Array of wires
assign mux[0] = input0; // Connects the sources of the array
assign mux[1] = input1;
assign mux[2] = input2;
assign mux[3] = input3;
assign mux[4] = input4;
assign mux[5] = input5;
assign mux[6] = input6;
assign mux[7] = input7;
assign mux[8] = input8;
assign mux[9] = input9;
assign mux[10] = input10;
assign mux[11] = input11;
assign mux[12] = input12;
assign mux[13] = input13;
assign mux[14] = input14;
assign mux[15] = input15;
assign mux[16] = input16;
assign mux[17] = input17;
assign mux[18] = input18;
assign mux[19] = input19;
assign mux[20] = input20;
assign mux[21] = input21;
assign mux[22] = input22;
assign mux[23] = input23;
assign mux[24] = input24;
assign mux[25] = input25;
assign mux[26] = input26;
assign mux[27] = input27;
assign mux[28] = input28;
assign mux[29] = input29;
assign mux[30] = input30;
assign mux[31] = input31;
assign out=mux[address]; // Connects the output of the array
endmodule


module decoder1to32(out, enable, address);
output[31:0] out;
input enable;
input[4:0] address;
assign out = enable<<address; //left shifts the enable bit however many bits the address declares
endmodule

module regfile(ReadData1, // Contents of first register read  //WORKED WITH LINDSEY ON THIS ONE
 ReadData2, // Contents of second register read
 WriteData, // Contents to write to register
 ReadRegister1, // Address of first register to read 
 ReadRegister2, // Address of second register to read
 WriteRegister, // Address of register to write
 RegWrite, // Enable writing of register when High
 Clk); // Clock (Positive Edge Triggered)

output[31:0] ReadData1, ReadData2;
input[4:0] ReadRegister1, ReadRegister2; //addresses of the two registers
input[31:0] WriteData; //0 or 1
input[4:0] WriteRegister; //address of the write
input Regwrite, Clk;

wire[31:0] decoderout;
wire[31:0] register[31:0];

decoder1to32 decoder1(decoderout, Regwrite, WriteRegister);
generate //Use generate to create an xor gate to check every bit
genvar index;
for (index = 0; index<32; index = index + 1)
	begin: regen
		register32 reg32bit(register[index], WriteData, decoderout[index], clk);
	end
endgenerate


endmodule

module test;

reg d, wrenable, clk;
wire q;
register reg1test(q, d, wrenable, clk);
initial begin
$display("D  | ENABLE  |  CLK  |   Q  ");
clk=1;wrenable=1;d=1; #5000
$display("%b  |%b  |%b  |%b  ", d, wrenable, clk, q);
clk=1;wrenable=1;d=0; #5000
$display("%b  |%b  |%b  |%b  ", d, wrenable, clk, q);
clk=0;wrenable=1;d=1; #5000
$display("%b  |%b  |%b  |%b  ", d, wrenable, clk, q);
clk=1;wrenable=1;d=0; #5000
$display("%b  |%b  |%b  |%b  ", d, wrenable, clk, q);
clk=0;wrenable=1;d=1; #5000
$display("%b  |%b  |%b  |%b  ", d, wrenable, clk, q);
end
endmodule

module test32;
reg[31:0] d;
reg wrenable;
reg clk;
wire[31:0] q;

register32 reg32bittest(q, d, wrenable, clk);

initial begin
$display("Testing AND");
$display("A                                 B                                |  Out                                 |Zero|  Expected");
clk=1;wrenable=1;d=32'b00000000000000000000000000000000; #10000 //all 0's test
$display("%b  %b |  %b    | %b  |  00000000000000000000000000000000", clk, wrenable, d, q);
clk=0;wrenable=1;d=32'b11111111111111111111111111111111; #10000 //all 0's test
$display("%b  %b |  %b    | %b  |  00000000000000000000000000000000", clk, wrenable, d, q);
clk=1;wrenable=1;d=32'b00000000000000000000111111111111; #10000 //all 0's test
$display("%b  %b |  %b    | %b  |  00000000000000000000000000000000", clk, wrenable, d, q);
end

endmodule